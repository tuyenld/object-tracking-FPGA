library verilog;
use verilog.vl_types.all;
entity filter_medium_vlg_tst is
end filter_medium_vlg_tst;
