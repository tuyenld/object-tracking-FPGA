library verilog;
use verilog.vl_types.all;
entity edge_detec_vlg_tst is
end edge_detec_vlg_tst;
