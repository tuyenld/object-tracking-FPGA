library verilog;
use verilog.vl_types.all;
entity test_clk_tb is
end test_clk_tb;
